library ieee;
use ieee.std_logic_1164.all;
 
entity Systolic_Array_Matrix_Multiplication is
end Systolic_Array_Matrix_Multiplication;

architecture Systolic_Array_Matrix_Multiplication_arch of Systolic_Array_Matrix_Multiplication is

begin


end Systolic_Array_Matrix_Multiplication_arch;