library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Input_data_controller is
	port(	data_in: in STD_LOGIC_VECTOR(3 downto 0);
			data_ready : in STD_LOGIC);
end Input_data_controller;

architecture Input_data_controller_arch of Input_data_controller is

begin


end Input_data_controller_arch;

