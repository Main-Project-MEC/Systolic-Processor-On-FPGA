library IEEE;
use IEEE.STD_LOGIC_1164.all;

package mem_content is

-- content of m_0_0
constant m_0_0_0 : BIT_VECTOR := X"9A94D4AD3DA5B5B3494A5E7F5F52F4B7E85E86F55BD2599BBED556D0FA186008";
constant m_0_0_1 : BIT_VECTOR := X"00000012FD4A9064A212F0B44569BF76453534FFD37B9A99B5352DA9A945352A";
constant m_0_0_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_0_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_1
constant m_0_1_0 : BIT_VECTOR := X"8CEDE77380EE7714C866432D57265582E6CAA054C9540EDCCD2B6B37844E6B08";
constant m_0_1_1 : BIT_VECTOR := X"0000007C3995A229037D7FCEF399199AEB19D542318B68EAB319C098CE1319D9";
constant m_0_1_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_1_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_2
constant m_0_2_0 : BIT_VECTOR := X"92F586973F82F429A96D4F64537EC5C66DD8B8C5EB151DE87C895C36445C4718";
constant m_0_2_1 : BIT_VECTOR := X"00000052C44FD2B4A712EC5ED8BDD4FA5525FB9252615AFC9525F9492FC525FA";
constant m_0_2_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_2_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_3
constant m_0_3_0 : BIT_VECTOR := X"C0E5B63BFF2769008C646709642017108602F210D05C4C60E88C4C26454D0B9B";
constant m_0_3_1 : BIT_VECTOR := X"0000005092DDB23DD35198EFC1DB01DF6181DA02181648EC9181C80C0E6181C8";
constant m_0_3_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_3_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_4
constant m_0_4_0 : BIT_VECTOR := X"C0E5B711C00228848C646100633007006600E00CD01E8640628C0C8350670813";
constant m_0_4_1 : BIT_VECTOR := X"0000002C60000200446C0C45C08B90C76181DA0A180400EC9181CC0C0E5181C8";
constant m_0_4_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_4_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_5
constant m_0_5_0 : BIT_VECTOR := X"1220A1207F2409A149124C89655696B4E852C29D5A5AD202A250542545230551";
constant m_0_5_1 : BIT_VECTOR := X"00000041000407007FC014834506854D04244299424092240424452122042442";
constant m_0_5_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_5_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_6
constant m_0_6_0 : BIT_VECTOR := X"DA868408C001183549524880634486242890C485421A102A0494100001290119";
constant m_0_6_1 : BIT_VECTOR := X"0000003EFF03C0F0773E04234446040405B508D25B6C9284D5B509ADA855B50A";
constant m_0_6_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_6_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_0_7
constant m_0_7_0 : BIT_VECTOR := X"00228000C000180048024000611006802200D004001800000240000001210011";
constant m_0_7_1 : BIT_VECTOR := X"0000000000000000000004034006800520004009000000204000400002000040";
constant m_0_7_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_0_7_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_0
constant m_1_0_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_1
constant m_1_1_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_2
constant m_1_2_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_3
constant m_1_3_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_4
constant m_1_4_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_5
constant m_1_5_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_6
constant m_1_6_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_7
constant m_1_7_0 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_1 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_2 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_3 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_8 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";


end mem_content;

package body mem_content is

end mem_content;

