library IEEE;
use IEEE.STD_LOGIC_1164.all;

package mem_content is

-- content of m_0_0
constant m_0_0_0 : BIT_VECTOR := X"E2BF124C93051303CFCCAC2652AEC692651B64AB6F4B926C081C0804080004D8";
constant m_0_0_1 : BIT_VECTOR := X"3FECF52100000231E7622B29268922F7931543E3664B3853387CEE7E65615B26";
constant m_0_0_2 : BIT_VECTOR := X"A3DF7793B9EFA732AAA25225224A0504A18029D278325DA4C200000709A03C38";
constant m_0_0_3 : BIT_VECTOR := X"16FB6E31C79C5674A32FF38CBCDDCC3AC9249D44A8BC952CC48B890935196A2A";
constant m_0_0_4 : BIT_VECTOR := X"9747FF77CA23FDFFD5BFFD5AA5FFEAD447FFAB5019BBED52FFDD5F2099A8D485";
constant m_0_0_5 : BIT_VECTOR := X"BEBDD5F1A999ABDED9BDB7E3C3C87F7FECF6FFECF7BDB97FF67BDED8BFFB3DEF";
constant m_0_0_6 : BIT_VECTOR := X"F5795E5795A769DE72DEF5AFDAA92E593BEBF001E1A9DD5E15659B6EFA4B6B57";
constant m_0_0_7 : BIT_VECTOR := X"C979FFA375642725E137AB37725E7FE8DD5909287E2725E7FECDD49094D55FD7";
constant m_0_0_8 : BIT_VECTOR := X"CC29BD98577B30A6F6615DECC5056F6418B3E6AF158EE4EE2725E7FE8DD49096";
constant m_0_0_9 : BIT_VECTOR := X"A9468AB07F9A8DD52A43627DAB64EFEB6142615DECC29BD98577B30A6F6615DE";
constant m_0_0_A : BIT_VECTOR := X"C37F407497FFC07C6F39FD9ABA7747C65D0AB43A1468556A56BA4AF04870D26E";
constant m_0_0_B : BIT_VECTOR := X"D5A1521A956A49666EFB555B43EA964B4EA54B4A2940E47252C115963FB6E0D3";
constant m_0_0_C : BIT_VECTOR := X"D914D4D3FF4DEE6A66D4D4B6A6A514D4AA6A5352B4F696CACD252979E92D4A92";
constant m_0_0_D : BIT_VECTOR := X"FB783C1E0F07825B7DA5A8B56DFEB66D412888104BF52A4192884BC2D115A6FD";
constant m_0_0_E : BIT_VECTOR := X"D949482400AE5242865241948065201242A2A48250A884F290DF6942A59554A6";
constant m_0_0_F : BIT_VECTOR := X"E37FFEB6A42ADBBBB776EDDCABFC921BF5B5247F1241E46A40934A52921525BE";

-- content of m_0_1
constant m_0_1_0 : BIT_VECTOR := X"80710228CA648A1C4AC88A359072F4E3512A2443C653894400000400080005F8";
constant m_0_1_1 : BIT_VECTOR := X"2CDA76114000020319D9E2815261D81190833D5B640CA648A1C4A25E44519435";
constant m_0_1_2 : BIT_VECTOR := X"584711D108232251871523DA353AE97B250035ADC4767BADF1000005A216E21B";
constant m_0_1_3 : BIT_VECTOR := X"227805D04096659DA10D7682C82A834F48844968961CC087A661488CA5A921C7";
constant m_0_1_4 : BIT_VECTOR := X"9050A52548A93452D3052D320429699010A5A64449CAD232525737A0D57AFD47";
constant m_0_1_5 : BIT_VECTOR := X"AF3C7AC2F0A8C7203045C2290F304D14A6AA14A6AB2A8B0A535594448529AACA";
constant m_0_1_6 : BIT_VECTOR := X"EF694EF694EF295EF2F7FDAFA41022C42AF0C8000EF6C7AD2F13A802BD1890E0";
constant m_0_1_7 : BIT_VECTOR := X"6156F7D6D11BD9855C9BA46D1855BDF1B446F6279219855BDF1B4C4E486CF694";
constant m_0_1_8 : BIT_VECTOR := X"633522C66E458CDC8B19A9163426C8B0464D9A22FF7BB0ABD9855BDF1B4C4E4A";
constant m_0_1_9 : BIT_VECTOR := X"A4EE4A88CA560B349EA159FA54B0ABB499BD99A91633522C66E458CDC8B19A91";
constant m_0_1_A : BIT_VECTOR := X"88093E5F9081BE5F9F2CA1A53F15F2360FDF1F9FBF3F1F3E7EEF2788D45AB659";
constant m_0_1_B : BIT_VECTOR := X"0F9B3A81D327503B7334ADACDE1FC8E55E10E44B0CAE7331395EC7A39F805D7E";
constant m_0_1_C : BIT_VECTOR := X"6BAC675508C62DA3AACC670263384C676633B79DCE03B9D45321990CBD7C99D6";
constant m_0_1_D : BIT_VECTOR := X"26F47A3D1E8F472B1372BDCC034A00E323915631F0E65688A40DF5FF3BCE6466";
constant m_0_1_E : BIT_VECTOR := X"A944E733BE62199C6A39D88E746399D9984833392E4E6BE9CEC4DCAAB2230E56";
constant m_0_1_F : BIT_VECTOR := X"F49B5E4973A800AD5564D56C292E39D350019D254333583B3249792C4E1F9989";

-- content of m_0_2
constant m_0_2_0 : BIT_VECTOR := X"094339A22811E831226222911943600815C01222E322D910000000040FFFFAD8";
constant m_0_2_1 : BIT_VECTOR := X"8021119540000264311108A4D1D45A49D84AB11170E2851E8712291311144691";
constant m_0_2_2 : BIT_VECTOR := X"3D374DDCCE9BB99CF4C89A01A01246517C0028D20D0300221940000404400681";
constant m_0_2_3 : BIT_VECTOR := X"810CD0934E45111006D2F323B23B637CA7D346F226C3D1A0516CA6A28BC21314";
constant m_0_2_4 : BIT_VECTOR := X"0B8A117245658508C3508C357284618A8A1186AA2C85C8D8882CD34A228540D4";
constant m_0_2_5 : BIT_VECTOR := X"5943E85C8A2008F70B2E687C38E7E1422E41422E41905CA11720C92F508B9064";
constant m_0_2_6 : BIT_VECTOR := X"4212908421480090004B1283B5B966C925DE97FFF9D83E8540F220416447DC3C";
constant m_0_2_7 : BIT_VECTOR := X"49BDDA54D2B72126FB52A54D126F769534ADC8973A9126F769134BFDA8488400";
constant m_0_2_8 : BIT_VECTOR := X"309790612B20C2564184AC830C52E418E1E3061C321924972126F769134BFDAA";
constant m_0_2_9 : BIT_VECTOR := X"2216631A98006004406B91BB5124972684B204AC8309590612F20C25E4184BC8";
constant m_0_2_A : BIT_VECTOR := X"4A211611561106100323C842E00B1C5E1C78C138718250A30EB8101A0D440300";
constant m_0_2_B : BIT_VECTOR := X"19B762E317AC5477A1F22570D9185A2D04342D13D5AE2699AB1EEC0149842C44";
constant m_0_2_C : BIT_VECTOR := X"E95497EE4949856BF25497E524BF1497EA4BD61A5CFE0BD8A6A5B53D914DFB17";
constant m_0_2_D : BIT_VECTOR := X"F60D068341A0D168FB16349044226A2428B156294B113F4AD29C4BB17B62F753";
constant m_0_2_E : BIT_VECTOR := X"A54C2D563E732B5A730B5EC2C770B12B1A5A56396D4562385A3EC58AD6ABA2C1";
constant m_0_2_F : BIT_VECTOR := X"C36DEC041630105D0BAD42EE59AC8B5B4022B535156365F16B6D129184F0B07D";

-- content of m_0_3
constant m_0_3_0 : BIT_VECTOR := X"0006843D0F080F409E1D1E5F1004CFC4F5074E20000011F80C0C0C0C000000C9";
constant m_0_3_1 : BIT_VECTOR := X"0CD2700740000109524077C210821021C00020405E10F080F40BE4F0E8F23C5F";
constant m_0_3_2 : BIT_VECTOR := X"28A7A1C00043800020044044044B6099BF800892559008B04060000106602AD8";
constant m_0_3_3 : BIT_VECTOR := X"10204088A13C8F26D0807802802A03721D084001040001020840909080000200";
constant m_0_3_4 : BIT_VECTOR := X"6121110490004488BB088BB000445DA10111768402088800884442241140C459";
constant m_0_3_5 : BIT_VECTOR := X"88054C008C465A2200603120BA379122209C22209C270A11104E128008882709";
constant m_0_3_6 : BIT_VECTOR := X"31CC731CE67B8EF399A5215935B92A5BC88137FFF96054C00111404232488000";
constant m_0_3_7 : BIT_VECTOR := X"9ED7DB6CD5166A7B5112AECD67B5F6DB35459A569D0A7B5F6DB35559AD99B9CF";
constant m_0_3_8 : BIT_VECTOR := X"9654272CA84E59509CB2A13965CA89CB2DF9F2E990C84F226A7B5F6DF35559AD";
constant m_0_3_9 : BIT_VECTOR := X"B4E7828B938683369A2EF4934B4F2246B2A6B2B139656272CA84E59509CB2A13";
constant m_0_3_A : BIT_VECTOR := X"DA1165E7451175E613AC8806CE11212710C91321932642644FC4A6AB45983619";
constant m_0_3_B : BIT_VECTOR := X"4C1833C98346713183A231309912AD57EC2057C00AD8443015F089D098044A1D";
constant m_0_3_C : BIT_VECTOR := X"7D86076808605923B246072030398607230396D8EFFC9DB80231919C39E0819C";
constant m_0_3_D : BIT_VECTOR := X"BF75BA5D6EB74AB55FABCC984223222E0D5F7475424B76C8F74D4663BF076C07";
constant m_0_3_E : BIT_VECTOR := X"E0A856ABE24015F06015B0056C015B15F0606B65887252C8AF57EAFD2BEF357A";
constant m_0_3_F : BIT_VECTOR := X"64891C042B60108F9124647C0C8C95E840215B9192B645CEBE498A5292E55EAF";

-- content of m_0_4
constant m_0_4_0 : BIT_VECTOR := X"00848018060306401898780C00840DC0C0461C20800010CC180C080C07FFF811";
constant m_0_4_1 : BIT_VECTOR := X"4C814146000001000211460000800600E08000014C006430600180C4C3C0F00C";
constant m_0_4_2 : BIT_VECTOR := X"200380E09001C120298C92C92C9B24480300000001B2990284600000064000D8";
constant m_0_4_3 : BIT_VECTOR := X"10014208A0303C2200A07A48A08A5800B9000500618231604018800014010200";
constant m_0_4_4 : BIT_VECTOR := X"210050F1B09000282082820A2814105100504145000028448C00406132050118";
constant m_0_4_5 : BIT_VECTOR := X"04202449CC440810612531088000000A1E340A1E358D00050F1AC68002878D63";
constant m_0_4_6 : BIT_VECTOR := X"6B58C6B5AD210A42918D695B74CB6ECBC0419000000802449809414010404994";
constant m_0_4_7 : BIT_VECTOR := X"5E00493A0C40E97805060BA05780124E83103A12B409780124E83103A50A158C";
constant m_0_4_8 : BIT_VECTOR := X"82018D04031A080634100C682F406341048B568CB65B2F00E9780124A83103A7";
constant m_0_4_9 : BIT_VECTOR := X"2297422300865324508C8437492F0127900E900C682018D04031A080634100C6";
constant m_0_4_A : BIT_VECTOR := X"530050C04050D0C003A20C20020010971C48913811227160C722142311843099";
constant m_0_4_B : BIT_VECTOR := X"0D983381B3467A19018A30320D402513802C13A80270241004A0001003142001";
constant m_0_4_C : BIT_VECTOR := X"1D86076828601003B246073030394607230396DC470008B21231918419ECC19C";
constant m_0_4_D : BIT_VECTOR := X"19008040603018940489C60060A0A00A8C4A224CB18000080111B03117022E43";
constant m_0_4_E : BIT_VECTOR := X"44A81289C00404A60404A90128404E84A60609C0002000002501225509492128";
constant m_0_4_F : BIT_VECTOR := X"2008011409545002000400100A8084EE08A04E50909C040094009294A6004A06";

-- content of m_0_5
constant m_0_5_0 : BIT_VECTOR := X"528E81485241520A28282814528C94914452148AA94A42540400000407FFF855";
constant m_0_5_1 : BIT_VECTOR := X"220104224000010146514A28A2A8A28ACA944A531405201520A2814141405114";
constant m_0_5_2 : BIT_VECTOR := X"8A2B8ACA8515950A28AA90A90A9344953900089251A055269260000141092840";
constant m_0_5_3 : BIT_VECTOR := X"04A32A28A050146680A93A4225200232A822955428A29428428A8505155148A8";
constant m_0_5_4 : BIT_VECTOR := X"64344AF1D2AA082504225040A5128204144A08145028250425414244AA0D1419";
constant m_0_5_5 : BIT_VECTOR := X"82151128A1112288108484AA728F82095E34895E358D2944AF1AC791A2578D63";
constant m_0_5_6 : BIT_VECTOR := X"635AC6B1AD6B58C6B18C63084A201800282247FFF52151120504532A0A082042";
constant m_0_5_7 : BIT_VECTOR := X"014124892D04940506E11892C05049224B41250A4D2405049224B4125108B18D";
constant m_0_5_8 : BIT_VECTOR := X"880B8D10171A202E34405C68830163441020C1AA010080A09405049264B41251";
constant m_0_5_9 : BIT_VECTOR := X"020748A13210088042065284A000A0894049405C6880B8D10171A202E34405C6";
constant m_0_5_A : BIT_VECTOR := X"3142D144544A41442B0A250AC85042864552A51A840A3448970210A140908044";
constant m_0_5_B : BIT_VECTOR := X"D5A1530AB56A6B480A89415095128141808541AAA832A15250651944A0328295";
constant m_0_5_C : BIT_VECTOR := X"3410910A6509024890109114848810910848828481FC902A8524493229A55A9A";
constant m_0_5_D : BIT_VECTOR := X"9951A8D46A151A054CA04A212894952A4D0223450400101C01FF00520D141A15";
constant m_0_5_E : BIT_VECTOR := X"456140A0CAA15062815068541A1502102282A0CA52829482835328332040040A";
constant m_0_5_F : BIT_VECTOR := X"204110B2A042CA8610468435A2501062A595064A820CA1CA0492108424E502A6";

-- content of m_0_6
constant m_0_6_0 : BIT_VECTOR := X"516CAA4E935593534C4EADA6516C66DA641B46AA4E4A9A600000000407FFF859";
constant m_0_6_1 : BIT_VECTOR := X"0CEB6412000001484604134D284D2AD2D21B521366A935593534DA62756D59A6";
constant m_0_6_2 : BIT_VECTOR := X"B34BD2D289A5A51296ACC0CC0CDB709981800A52109A0892512000001660085C";
constant m_0_6_3 : BIT_VECTOR := X"16AA4A2AAA9B5662240D7A10800A00800DB49466AAA8D5AA54AA296941946B36";
constant m_0_6_4 : BIT_VECTOR := X"742692719A82AB496434964281A4B2140692C85412A049402901093011A49008";
constant m_0_6_5 : BIT_VECTOR := X"021015A82DDDA88A14B0B68340882AD24E36D24E378DA869271BC7D534938DE3";
constant m_0_6_6 : BIT_VECTOR := X"214A5210A5294A5231AC6B1D92ADAB61A02040000109015A84441A4808622042";
constant m_0_6_7 : BIT_VECTOR := X"0D012499244524340921499243404926491149A95514340492649114930A94A4";
constant m_0_6_8 : BIT_VECTOR := X"E8A98DD1531BA2A637454C6E8515637450A142A2110886812434049264911493";
constant m_0_6_9 : BIT_VECTOR := X"B6C74A2120974336D8040299200680824552454C6E8A98DD1531BA2A637454C6";
constant m_0_6_A : BIT_VECTOR := X"126A52611692D261232029A8004042065D52A52AA54A550A1700B6010080B819";
constant m_0_6_B : BIT_VECTOR := X"90A2431215086840A81250400000211184B511A32234A6514469501722A48484";
constant m_0_6_C : BIT_VECTOR := X"1016D423496DB24A1356D426B6A156D42B6A1A1023000468D5254922018D1218";
constant m_0_6_D : BIT_VECTOR := X"0B0080402010088C058842A14D25241A24426644FBFC0F03C1DCF8108D111810";
constant m_0_6_E : BIT_VECTOR := X"D16D1088D4A2446AA2446091182446046A8A885294ACA4022101623308CC3118";
constant m_0_6_F : BIT_VECTOR := X"2248842488C092028054A0102C94C42AA12442929884A60084921AD6B7004202";

-- content of m_0_7
constant m_0_7_0 : BIT_VECTOR := X"0080010842414248282829141080148141020400210040400000000400000241";
constant m_0_7_1 : BIT_VECTOR := X"0A8340020000000800150A208A208208C8840800140420142082914141485014";
constant m_0_7_2 : BIT_VECTOR := X"082388C804119008888210210203148401000240008804020020000015400054";
constant m_0_7_3 : BIT_VECTOR := X"0021220000521400008038400402400088020010208010200208044440400088";
constant m_0_7_4 : BIT_VECTOR := X"6020484010800224000240002012000100480000000024000400091008040108";
constant m_0_7_5 : BIT_VECTOR := X"0000000800000082041400200080008908040908040100048402008002420100";
constant m_0_7_6 : BIT_VECTOR := X"214A52948421084210A521084804892800081000040000000000012000200000";
constant m_0_7_7 : BIT_VECTOR := X"4010000804409100448048805004000201102400040100400020100241421084";
constant m_0_7_8 : BIT_VECTOR := X"8202010404020808041010082140004104085080804020009100400020100241";
constant m_0_7_9 : BIT_VECTOR := X"06874021008542A0D08410048920002910091010082020104040208080410100";
constant m_0_7_A : BIT_VECTOR := X"11005141004851410B0000020200109604000008000010000700342110802815";
constant m_0_7_B : BIT_VECTOR := X"04881340900260000009000000000300A0040080801201000024000080120204";
constant m_0_7_C : BIT_VECTOR := X"1480010024000000810001000008000100008A00030000680120090009A4409A";
constant m_0_7_D : BIT_VECTOR := X"090080402010080C0480C208209091100406664C00000000000000100D001A00";
constant m_0_7_E : BIT_VECTOR := X"406001804A210022210028400A10028022220048420210000101203300C82018";
constant m_0_7_F : BIT_VECTOR := X"2248801200D04802801020140244406200900648080C22000C00000001000602";

-- content of m_1_0
constant m_1_0_0 : BIT_VECTOR := X"E5E0924F05AD3BEC52829CFDAFFF7EFFAF2B5FD201E0900D20B7B41DE0924832";
constant m_1_0_1 : BIT_VECTOR := X"04A24A04964929EFCFD28E74A2E9673A5934F4A39D2CABA4B16D65E03F249241";
constant m_1_0_2 : BIT_VECTOR := X"8A412056D752A9E02F7BD752A9E02F73D09E0F04824124920C0E9E0944555535";
constant m_1_0_3 : BIT_VECTOR := X"000001E3C3777EAB7773F56EEC7BADDDCA9078241EA78249549176D5B5AA48A4";
constant m_1_0_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_8 : BIT_VECTOR := X"880140807C6807C6803A2C000000000000000000000000000000000000000000";
constant m_1_0_9 : BIT_VECTOR := X"801CE4B9C536A49F2B8E0029E91F562502C2982B550056AA53E19B235C46394F";
constant m_1_0_A : BIT_VECTOR := X"4895717C7129B6C4810133C1085B924C90C9A388000A2E3310AE4EA0AE239675";
constant m_1_0_B : BIT_VECTOR := X"5F47CD474F6ABF32B73D539E882248FB762D558A32E44D0BC944CC72B4B9571C";
constant m_1_0_C : BIT_VECTOR := X"E31C831C849DC891DC85115F2D5048D56322B9195BD5AB46ADECC8F355D5C2EE";
constant m_1_0_D : BIT_VECTOR := X"00000000000000000000000000000000000000000000000000000000724AC77C";
constant m_1_0_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_0_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_1
constant m_1_1_0 : BIT_VECTOR := X"931179D88A1ECA9082DEDFAD29DAD2BDE73BDB351F10CCEB5038631311CCD440";
constant m_1_1_1 : BIT_VECTOR := X"8E75677ACCF79C1D7439D3AE751CEDD732FB0E74EB98965E76CA305BF95E76A3";
constant m_1_1_2 : BIT_VECTOR := X"B6A351492202815BFC9F2AA6D35BFC972F31188E46A04135100EF11CCB2AAA84";
constant m_1_1_3 : BIT_VECTOR := X"0000017E215953EA557A7D4AAD4AA955A9A8C46A22DC432A0654255320A32A32";
constant m_1_1_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000100000";
constant m_1_1_8 : BIT_VECTOR := X"A8012080330804A680330E000000000000000000000000000000000000000000";
constant m_1_1_9 : BIT_VECTOR := X"4002C943DB0B492E3096001832E8624B8480A04C660098CC30608537586EB0C1";
constant m_1_1_A : BIT_VECTOR := X"1C296235629D20280E24574421100489948022940017300000309420C2110A65";
constant m_1_1_B : BIT_VECTOR := X"281B8D0AC168C81056346B1A310501494C08881022608086110808A034380628";
constant m_1_1_C : BIT_VECTOR := X"C12009200829420294112FA852B801220084980466090502130081034601826C";
constant m_1_1_D : BIT_VECTOR := X"00000000000000000000000000000000000000000000000000000000601988A0";
constant m_1_1_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_1_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_2
constant m_1_2_0 : BIT_VECTOR := X"78348B01A5C785C90F250000520425210042148348355AE034FD8E38345A0D3F";
constant m_1_2_1 : BIT_VECTOR := X"A2C2AD5558A8B4611C4B48E2D2258471691E12C238B1CBAAD4E48139EF22C068";
constant m_1_2_2 : BIT_VECTOR := X"B06834A086360939E3B0E6360939E3B0E08341A2E06B64834FFC8345A5575508";
constant m_1_2_3 : BIT_VECTOR := X"0000011068B0B9220B0204416040882C481A0D069F20D57ACAF4720392157357";
constant m_1_2_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000080000";
constant m_1_2_8 : BIT_VECTOR := X"88016000664807C6001F28000000000000000000000000000000000000000000";
constant m_1_2_9 : BIT_VECTOR := X"001A14B8F744A490B4BC0028C9FA6B2F864E18707800E0F051ABA26E02DC0546";
constant m_1_2_A : BIT_VECTOR := X"0DCC09C009E81544850F2E8F7BC35245A859C118001F167733964B40D2B69009";
constant m_1_2_B : BIT_VECTOR := X"53442C5546623A5A208110408863F0A6376165CA01424E83C8E42256899DF194";
constant m_1_2_C : BIT_VECTOR := X"159D859D871619E1618B9F9329D988D9752A50A913CBAAECA9E22AEB117C6141";
constant m_1_2_D : BIT_VECTOR := X"000000000000000000000000000000000000000000000000000000000B8DDF4C";
constant m_1_2_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_2_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_3
constant m_1_3_0 : BIT_VECTOR := X"155615EA90AC88E810208563085694842148C6112952AF9D12B0BB5152AD44CF";
constant m_1_3_1 : BIT_VECTOR := X"357856D0ADA15F117515ABA5788AF5D2B432456AE95EA2056C89515CA9057A2D";
constant m_1_3_2 : BIT_VECTOR := X"E22516808E995E5CA8922E995E5CA89220956A956A252D9133F2152AD1061028";
constant m_1_3_3 : BIT_VECTOR := X"00000052A51D1C621102AC42225188444A8955A2E5A54AB7456C44EA2542B62B";
constant m_1_3_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_8 : BIT_VECTOR := X"D00141002E3800D3806552000000000000000000000000000000000000000000";
constant m_1_3_9 : BIT_VECTOR := X"800A8DE26151EDB41A14000C9BE3336B86001201800403001930A86610CC2064";
constant m_1_3_A : BIT_VECTOR := X"0848432C4388860C94346614A50986C198404010001704004004D80068500C41";
constant m_1_3_B : BIT_VECTOR := X"014D064C6432631AE42D3216995715940004011D1484C20B582CA4C098388834";
constant m_1_3_C : BIT_VECTOR := X"81B009B00AB2822B28193EC17C14AB80402721013B55AE209DAA49B193A21488";
constant m_1_3_D : BIT_VECTOR := X"00000000000000000000000000000000000000000000000000000000414BCA04";
constant m_1_3_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_3_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_4
constant m_1_4_0 : BIT_VECTOR := X"044304E218A00029326DEE399EF398C73BDE72047046251847B8885046251180";
constant m_1_4_1 : BIT_VECTOR := X"312C128827104A801084A8813C4270409E00213A204AB1412863C18208412884";
constant m_1_4_2 : BIT_VECTOR := X"408C438287188C82000007188C82000008842231288D2484200104627820823A";
constant m_1_4_3 : BIT_VECTOR := X"000000308C0407620022EC40045988008E23108840611895413871918D209409";
constant m_1_4_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_5 : BIT_VECTOR := X"0000000000000000000000000000000040000000000000000000000000000000";
constant m_1_4_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000180000";
constant m_1_4_8 : BIT_VECTOR := X"F0016180757807C5005F56000000000000000000000000000000000000000000";
constant m_1_4_9 : BIT_VECTOR := X"600050138A0A000A84A80012200000002484E301FF8603FF247B05184A309491";
constant m_1_4_A : BIT_VECTOR := X"D0012801281122201A3A105AD69070080082278C000038226138076012C18A0C";
constant m_1_4_B : BIT_VECTOR := X"3802A9129148800012804940218020684808EA45A168048C01009830A0044209";
constant m_1_4_C : BIT_VECTOR := X"50000800080882408812803802A1003A90885A044C10010A0609800A40108165";
constant m_1_4_D : BIT_VECTOR := X"00000000000000000000000000000000000000000000000000000000281410E0";
constant m_1_4_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_4_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_5
constant m_1_5_0 : BIT_VECTOR := X"0D46902A346828214480842958C6B18C6B1A525069468129063221C54681418F";
constant m_1_5_1 : BIT_VECTOR := X"340A419481290282409022041A4835020D20A4188106682409635490A1241A0D";
constant m_1_5_2 : BIT_VECTOR := X"CA0D06B652422190A81202422190A81204146A341A0C001063F2146814924929";
constant m_1_5_3 : BIT_VECTOR := X"000000428D0505495041812A0A112541068351A0C4A51A0CD40931858F0A04A0";
constant m_1_5_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000080000";
constant m_1_5_8 : BIT_VECTOR := X"6804000029280090802228000000000000000000000000000000000000000000";
constant m_1_5_9 : BIT_VECTOR := X"DFFFE01FFEFC000FFF7DFFFFC0FFFE0FAFDFFB7FFF8203FF7FDBFF7FFEFFFDFF";
constant m_1_5_A : BIT_VECTOR := X"FFFFF0FFF0FFF001CFAF1FEF7BFFE01FC1FC0821FFFF7EFFBFFE07DFFFEF7DFB";
constant m_1_5_B : BIT_VECTOR := X"FFF3FFE3FFFF1FFF1FFFCFFFE7E1F87EFFFFFF83FFF01F5F8301FC3FE3FFFF8F";
constant m_1_5_C : BIT_VECTOR := X"EF0FFF8FFF8FFFF8FFFF8FFE07FE1C7FFFF9FC7FCFFFF91FE7FFFE7FFCFFFFFF";
constant m_1_5_D : BIT_VECTOR := X"00000000000000000000000000000000000000000000000000000000779F9FF9";
constant m_1_5_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_5_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_6
constant m_1_6_0 : BIT_VECTOR := X"4C02046010E2202954818C6B5AC6B5AC694843402002234C02B289D4022300A0";
constant m_1_6_1 : BIT_VECTOR := X"910811802300462A02046811080210088408810A0442E0010963650208811804";
constant m_1_6_2 : BIT_VECTOR := X"480402A4965AAD020248965AAD02024894C020110805B6C02800002210000828";
constant m_1_6_3 : BIT_VECTOR := X"000000100404044A40538948087029010A0100805000088DD11971958FA88C88";
constant m_1_6_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_8 : BIT_VECTOR := X"E80000802820008000020A000000000000000000000000000000000000000000";
constant m_1_6_9 : BIT_VECTOR := X"E01EF011FF7E000FBFBE003FE01F7F078088827E0004FC007FFBBF7F1EFE3DFF";
constant m_1_6_A : BIT_VECTOR := X"1DFC78FC787DA3E010101FD0841BF009BCD3E79C000F2044422007E0FEF79E7D";
constant m_1_6_B : BIT_VECTOR := X"7F13EF13FF789F7887BC03DE00F0FC7F7F4DFFC537EE0F8FC1E0FE343D3DFF8C";
constant m_1_6_C : BIT_VECTOR := X"F7810781078FD1F8FD0F81FF03F9E27FF789FBBC4FDF89EE27EFE27BC47FE7EF";
constant m_1_6_D : BIT_VECTOR := X"000000000000000000000000000000000000000000000000000000007BDFDFFC";
constant m_1_6_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_6_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";

-- content of m_1_7
constant m_1_7_0 : BIT_VECTOR := X"4442006210200021100084294A521084294A52042042032842300940420310A0";
constant m_1_7_1 : BIT_VECTOR := X"1018008001000280128020900840104804002008240220000800500008801884";
constant m_1_7_2 : BIT_VECTOR := X"C084420242000000024892000000024894442210188492442800042030020008";
constant m_1_7_3 : BIT_VECTOR := X"00000000840405010010A02002140400422110885001080C4018000001000C00";
constant m_1_7_4 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_5 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_6 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_7 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_8 : BIT_VECTOR := X"0805808008080000802228000000000000000000000000000000000000000000";
constant m_1_7_9 : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_A : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_B : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_C : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_D : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_E : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";
constant m_1_7_F : BIT_VECTOR := X"0000000000000000000000000000000000000000000000000000000000000000";


end mem_content;

package body mem_content is

end mem_content;

